* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : tristatebuffer_x1                            *
* Netlisted  : Tue Nov 25 20:16:17 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764112572790                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764112572790 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.46017 scb=0.000436376 scc=1.63659e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764112572790

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv_x1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv_x1 Vin Vout vdd! gnd!
** N=4 EP=4 FDC=2
X2 gnd! Vout Vin nmos1v_CDNS_764112572790 $T=640 820 0 0 $X=220 $Y=620
M0 Vout Vin vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=31.4202 scb=0.0358526 scc=0.00253079 $X=640 $Y=2850 $dt=1
.ends inv_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764112572792                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764112572792 1 2 3
** N=4 EP=3 FDC=1
M0 3 2 1 1 g45p1svt L=4.5e-08 W=1.45e-07 AD=8.7e-15 AS=2.03e-14 PD=4.1e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=2.45e-07 sca=26.5414 scb=0.0263556 scc=0.002507 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764112572792

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764112572793                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764112572793 1 2 3 5
** N=5 EP=4 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=8.7e-15 PD=5.7e-07 PS=4.1e-07 fw=1.45e-07 sa=2.45e-07 sb=1.4e-07 sca=27.3953 scb=0.0274124 scc=0.00251189 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764112572793

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764112572794                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764112572794 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=4.46017 scb=0.000436376 scc=1.63659e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764112572794

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764112572795                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764112572795 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=4.46017 scb=0.000436376 scc=1.63659e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764112572795

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: tristatebuffer_x1                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt tristatebuffer_x1 en gnd! in out vdd!
** N=9 EP=5 FDC=8
X5 gnd! 2 in nmos1v_CDNS_764112572790 $T=2200 820 0 0 $X=1780 $Y=620
X7 en 3 vdd! gnd! inv_x1 $T=0 0 0 0 $X=0 $Y=0
X8 vdd! 2 7 pmos1v_CDNS_764112572792 $T=3390 2830 0 0 $X=2970 $Y=2630
X9 out 3 7 vdd! pmos1v_CDNS_764112572793 $T=3600 2830 0 0 $X=3400 $Y=2630
X10 out en 9 gnd! nmos1v_CDNS_764112572794 $T=3600 820 0 0 $X=3400 $Y=620
X11 gnd! 2 9 nmos1v_CDNS_764112572795 $T=3390 820 0 0 $X=2970 $Y=620
M0 2 in vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=24.5515 scb=0.0251693 scc=0.00232652 $X=2200 $Y=2840 $dt=1
.ends tristatebuffer_x1

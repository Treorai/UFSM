* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : flipflopD_x1                                 *
* Netlisted  : Tue Nov 25 20:55:16 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_764114911960                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_764114911960 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_764114911960

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_764114911961                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_764114911961 1 2
** N=2 EP=2 FDC=0
.ends M1_NWELL_CDNS_764114911961

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764114911962                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764114911962 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764114911962

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764114911963                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764114911963 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764114911963

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764114911964                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764114911964 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764114911964

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764114911966                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764114911966 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764114911966

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764114911967                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764114911967 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764114911967

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764114911968                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764114911968 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764114911968

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764114911969                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764114911969 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764114911969

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764114911960                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764114911960 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.92313 scb=0.000827672 scc=8.57018e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764114911960

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764114911961                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764114911961 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_764114911961

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764114911962                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764114911962 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 3 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.32e-14 PD=5.7e-07 PS=6.1e-07 fw=1.45e-07 sa=3.45e-07 sb=1.4e-07 sca=22.508 scb=0.0238066 scc=0.00185903 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764114911962

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764114911963                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764114911963 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 3 1 1 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.32e-14 AS=2.03e-14 PD=6.1e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=3.45e-07 sca=22.508 scb=0.0238066 scc=0.00185903 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764114911963

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764114911964                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764114911964 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.32e-14 PD=5.7e-07 PS=6.1e-07 fw=1.45e-07 sa=3.45e-07 sb=1.4e-07 sca=22.508 scb=0.0238066 scc=0.00185903 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764114911964

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764114911965                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764114911965 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 3 1 1 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.32e-14 PD=5.7e-07 PS=6.1e-07 fw=1.45e-07 sa=3.45e-07 sb=1.4e-07 sca=22.508 scb=0.0238066 scc=0.00185903 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764114911965

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764114911966                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764114911966 1 2 3
** N=3 EP=3 FDC=1
M0 1 2 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=4.92313 scb=0.000827672 scc=8.57018e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764114911966

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764114911967                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764114911967 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=4.92313 scb=0.000827672 scc=8.57018e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764114911967

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: flipflopD_x1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt flipflopD_x1 9 8 10 4 1 2
** N=10 EP=6 FDC=12
X0 1 M1_PSUB_CDNS_764114911960 $T=4310 300 0 0 $X=1890 $Y=160
X1 2 1 M1_NWELL_CDNS_764114911961 $T=4300 3700 0 0 $X=1840 $Y=3400
X2 3 M1_PO_CDNS_764114911962 $T=1150 2380 0 90 $X=1030 $Y=2280
X3 4 M1_PO_CDNS_764114911962 $T=5150 1750 0 0 $X=5050 $Y=1630
X4 5 M1_PO_CDNS_764114911963 $T=1660 1590 0 0 $X=1320 $Y=1470
X5 6 M1_PO_CDNS_764114911963 $T=5240 2360 0 0 $X=4900 $Y=2240
X6 7 M2_M1_CDNS_764114911964 $T=2470 2150 0 0 $X=2250 $Y=2020
X7 6 M2_M1_CDNS_764114911964 $T=3320 2360 0 0 $X=3100 $Y=2230
X8 6 M2_M1_CDNS_764114911964 $T=5240 2360 0 0 $X=5020 $Y=2230
X9 4 M2_M1_CDNS_764114911964 $T=7930 2210 0 0 $X=7710 $Y=2080
X10 5 M2_M1_CDNS_764114911966 $T=1660 1590 0 0 $X=1300 $Y=1460
X11 8 M2_M1_CDNS_764114911966 $T=6940 2350 0 0 $X=6580 $Y=2220
X12 7 M2_M1_CDNS_764114911967 $T=4770 1760 0 180 $X=4690 $Y=1630
X13 6 M2_M1_CDNS_764114911967 $T=8040 1640 0 0 $X=7960 $Y=1510
X14 7 M3_M2_CDNS_764114911968 $T=2330 2150 0 0 $X=2250 $Y=2020
X15 7 M3_M2_CDNS_764114911968 $T=4770 1760 0 0 $X=4690 $Y=1630
X16 5 M2_M1_CDNS_764114911969 $T=3410 1270 0 0 $X=3330 $Y=1000
X17 4 M2_M1_CDNS_764114911969 $T=5150 1760 0 0 $X=5070 $Y=1490
X18 1 5 3 1 nmos1v_CDNS_764114911960 $T=720 1000 0 0 $X=300 $Y=800
X19 1 3 7 1 nmos1v_CDNS_764114911960 $T=2500 1000 0 0 $X=2080 $Y=800
X20 5 4 9 1 nmos1v_CDNS_764114911960 $T=4380 1000 0 0 $X=3960 $Y=800
X21 8 4 6 1 nmos1v_CDNS_764114911960 $T=7790 1000 0 0 $X=7370 $Y=800
X22 2 3 5 1 2 pmos1v_CDNS_764114911961 $T=720 2870 0 0 $X=300 $Y=2670
X23 5 7 4 1 2 pmos1v_CDNS_764114911961 $T=4380 2870 0 0 $X=3960 $Y=2670
X24 8 10 2 1 pmos1v_CDNS_764114911962 $T=6390 2870 0 0 $X=6150 $Y=2670
X25 2 7 3 1 pmos1v_CDNS_764114911963 $T=2500 2870 0 0 $X=2080 $Y=2670
X26 6 4 7 1 2 pmos1v_CDNS_764114911964 $T=2910 2870 0 0 $X=2670 $Y=2670
X27 2 10 6 1 pmos1v_CDNS_764114911965 $T=6070 2870 1 180 $X=5560 $Y=2670
X28 8 10 1 nmos1v_CDNS_764114911966 $T=6390 1000 0 0 $X=6150 $Y=800
X29 1 10 6 nmos1v_CDNS_764114911967 $T=6070 1000 1 180 $X=5560 $Y=800
M0 3 5 2 2 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=28.4097 scb=0.0321484 scc=0.00204568 $X=720 $Y=2870 $dt=1
M1 7 4 5 2 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=22.508 scb=0.0238066 scc=0.00185903 $X=4380 $Y=2870 $dt=1
.ends flipflopD_x1

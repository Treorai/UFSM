************************************************************************
* auCdl Netlist:
* 
* Library Name:  watto
* Top Cell Name: 1_bit_full_adder_x1
* View Name:     schematic
* Netlisted on:  Dec  1 22:52:56 2025
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL vdd!
+        gnd!

*.PIN vdd!
*+    gnd!

************************************************************************
* Library Name: watto
* Cell Name:    nand_x1
* View Name:    schematic
************************************************************************

.SUBCKT nand_x1 A B S
*.PININFO A:I B:I S:O
MPM1 vdd! B S vdd! g45p1svt m=1 l=45n w=145n
MPM0 S A vdd! vdd! g45p1svt m=1 l=45n w=145n
MNM1 net9 B gnd! gnd! g45n1svt m=1 l=45n w=120n
MNM0 S A net9 gnd! g45n1svt m=1 l=45n w=120n
.ENDS

************************************************************************
* Library Name: watto
* Cell Name:    1_bit_full_adder_x1
* View Name:    schematic
************************************************************************

.SUBCKT 1_bit_full_adder_x1 A B CarryIn CarryOut S
*.PININFO A:I B:I CarryIn:I CarryOut:O S:O
XI8 net15 net3 CarryOut / nand_x1
XI7 net18 net21 S / nand_x1
XI6 net15 CarryIn net21 / nand_x1
XI5 net12 net15 net18 / nand_x1
XI4 net12 CarryIn net15 / nand_x1
XI3 net6 net9 net12 / nand_x1
XI2 net3 B net9 / nand_x1
XI1 A net3 net6 / nand_x1
XI0 A B net3 / nand_x1
.ENDS


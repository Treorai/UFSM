* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : 1_bit_full_adder_x1                          *
* Netlisted  : Mon Dec  1 22:53:01 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764640374440                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764640374440 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 3 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.74923 scb=0.000663449 scc=4.92991e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764640374440

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nand_x1                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nand_x1 B A S vdd! gnd!
*.DEVICECLIMB
** N=6 EP=5 FDC=2
X9 gnd! 6 B gnd! nmos1v_CDNS_764640374440 $T=860 940 0 0 $X=440 $Y=740
X10 6 S A gnd! nmos1v_CDNS_764640374440 $T=2260 940 0 0 $X=1840 $Y=740
.ends nand_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 1_bit_full_adder_x1                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 1_bit_full_adder_x1 A B CarryIn CarryOut S gnd! vdd!
** N=23 EP=7 FDC=36
X17 B A 2 vdd! gnd! nand_x1 $T=0 0 0 0 $X=0 $Y=0
X18 B 2 9 vdd! gnd! nand_x1 $T=3210 0 0 0 $X=3210 $Y=0
X19 9 3 4 vdd! gnd! nand_x1 $T=6420 0 0 0 $X=6420 $Y=0
X20 2 A 3 vdd! gnd! nand_x1 $T=9630 0 0 0 $X=9630 $Y=0
X21 CarryIn 4 11 vdd! gnd! nand_x1 $T=12840 0 0 0 $X=12840 $Y=0
X22 CarryIn 11 5 vdd! gnd! nand_x1 $T=16050 0 0 0 $X=16050 $Y=0
X23 2 11 CarryOut vdd! gnd! nand_x1 $T=19260 0 0 0 $X=19260 $Y=0
X24 11 4 13 vdd! gnd! nand_x1 $T=22470 0 0 0 $X=22470 $Y=0
X25 5 13 S vdd! gnd! nand_x1 $T=25680 0 0 0 $X=25680 $Y=0
M0 2 A vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=33.2274 scb=0.0325337 scc=0.00341592 $X=860 $Y=2790 $dt=1
M1 vdd! B 2 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=2260 $Y=2790 $dt=1
M2 9 2 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=4070 $Y=2790 $dt=1
M3 vdd! B 9 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=5470 $Y=2790 $dt=1
M4 4 3 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=7280 $Y=2790 $dt=1
M5 vdd! 9 4 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=8680 $Y=2790 $dt=1
M6 3 A vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=10490 $Y=2790 $dt=1
M7 vdd! 2 3 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=11890 $Y=2790 $dt=1
M8 11 4 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=13700 $Y=2790 $dt=1
M9 vdd! CarryIn 11 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=15100 $Y=2790 $dt=1
M10 5 11 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=16910 $Y=2790 $dt=1
M11 vdd! CarryIn 5 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=18310 $Y=2790 $dt=1
M12 CarryOut 11 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=20120 $Y=2790 $dt=1
M13 vdd! 2 CarryOut vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=21520 $Y=2790 $dt=1
M14 13 4 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=23330 $Y=2790 $dt=1
M15 vdd! 11 13 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=24730 $Y=2790 $dt=1
M16 S 13 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.2883 scb=0.0276453 scc=0.0033614 $X=26540 $Y=2790 $dt=1
M17 vdd! 5 S vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=33.2274 scb=0.0325337 scc=0.00341592 $X=27940 $Y=2790 $dt=1
.ends 1_bit_full_adder_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : flipflopD_x1                                 *
* Netlisted  : Mon Dec  1 16:49:26 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764618561424                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764618561424 1 2 3 5
** N=5 EP=4 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=8.7e-15 PD=5.7e-07 PS=4.1e-07 fw=1.45e-07 sa=2.45e-07 sb=1.4e-07 sca=25.5193 scb=0.0270883 scc=0.00188132 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764618561424

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764618561425                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764618561425 1 2 3
** N=4 EP=3 FDC=1
M0 3 2 1 1 g45p1svt L=4.5e-08 W=1.45e-07 AD=8.7e-15 AS=2.03e-14 PD=4.1e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=2.45e-07 sca=27.9002 scb=0.0312654 scc=0.00200277 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764618561425

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764618561426                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764618561426 1 2 3
** N=4 EP=3 FDC=1
M0 3 2 1 1 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.32e-14 AS=2.03e-14 PD=6.1e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=3.45e-07 sca=22.508 scb=0.0238066 scc=0.00185903 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764618561426

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764618561427                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764618561427 1 2 3
** N=4 EP=3 FDC=1
M0 1 3 2 2 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.32e-14 AS=2.03e-14 PD=6.1e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=3.45e-07 sca=22.508 scb=0.0238066 scc=0.00185903 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764618561427

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: flipflopD_x1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt flipflopD_x1 D Q Reset clk gnd! vdd!
** N=12 EP=6 FDC=12
X13 9 clk 12 vdd! pmos1v_CDNS_764618561424 $T=960 2870 0 0 $X=760 $Y=2670
X14 vdd! D 12 pmos1v_CDNS_764618561425 $T=750 2870 0 0 $X=330 $Y=2670
X15 vdd! Reset 5 pmos1v_CDNS_764618561426 $T=4370 2870 1 180 $X=4040 $Y=2670
X16 5 vdd! 6 pmos1v_CDNS_764618561427 $T=3870 2870 0 0 $X=3450 $Y=2670
M0 9 D gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=5.43278 scb=0.00141223 scc=3.10179e-06 $X=750 $Y=1140 $dt=0
M1 10 clk gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=5.34932 scb=0.00130706 scc=2.58259e-06 $X=2680 $Y=1120 $dt=0
M2 6 9 10 gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=5.34932 scb=0.00130706 scc=2.58259e-06 $X=2890 $Y=1120 $dt=0
M3 11 clk 5 gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=5.30908 scb=0.00125757 scc=2.35636e-06 $X=4280 $Y=1110 $dt=0
M4 gnd! 6 11 gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=5.30908 scb=0.00125757 scc=2.35636e-06 $X=4490 $Y=1110 $dt=0
M5 Q 5 gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=5.30908 scb=0.00125757 scc=2.35636e-06 $X=5800 $Y=1110 $dt=0
M6 6 clk vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=23.1359 scb=0.0242481 scc=0.00200358 $X=2360 $Y=2860 $dt=1
M7 Q 5 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.3403 scb=0.0285068 scc=0.00190891 $X=5800 $Y=2870 $dt=1
.ends flipflopD_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : buffer_x2                                    *
* Netlisted  : Tue Nov 25 18:37:27 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764106643070                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764106643070 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=4.82293 scb=0.000845673 scc=1.19259e-06 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764106643070

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764106643071                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764106643071 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_764106643071

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv_x2                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv_x2 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X0 4 2 1 nmos1v_CDNS_764106643070 $T=640 820 0 0 $X=220 $Y=620
X1 3 2 1 4 pmos1v_CDNS_764106643071 $T=640 2580 0 0 $X=220 $Y=2380
.ends inv_x2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: buffer_x2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt buffer_x2 4 1 5 3
** N=5 EP=4 FDC=4
X0 1 2 3 4 inv_x2 $T=0 0 0 0 $X=0 $Y=0
X1 2 5 3 4 inv_x2 $T=1550 0 0 0 $X=1550 $Y=0
M0 2 1 3 3 g45p1svt L=4.5e-08 W=2.9e-07 AD=4.06e-14 AS=4.06e-14 PD=8.6e-07 PS=8.6e-07 fw=2.9e-07 sa=1.4e-07 sb=1.4e-07 sca=60.4911 scb=0.0392764 scc=0.00603914 $X=640 $Y=2580 $dt=1
M1 5 2 3 3 g45p1svt L=4.5e-08 W=2.9e-07 AD=4.06e-14 AS=4.06e-14 PD=8.6e-07 PS=8.6e-07 fw=2.9e-07 sa=1.4e-07 sb=1.4e-07 sca=61.0162 scb=0.0400902 scc=0.00610802 $X=2190 $Y=2580 $dt=1
.ends buffer_x2

************************************************************************
* auCdl Netlist:
* 
* Library Name:  watto
* Top Cell Name: nor_x1
* View Name:     schematic
* Netlisted on:  Nov 26 23:24:32 2025
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL vdd!
+        gnd!

*.PIN vdd!
*+    gnd!

************************************************************************
* Library Name: watto
* Cell Name:    nor_x1
* View Name:    schematic
************************************************************************

.SUBCKT nor_x1 A B S
*.PININFO A:I B:I S:O
MPM1 net6 A S vdd! g45p1svt m=1 l=45n w=145n
MPM0 net6 B vdd! vdd! g45p1svt m=1 l=45n w=145n
MNM1 S B gnd! gnd! g45n1svt m=1 l=45n w=120n
MNM0 S A gnd! gnd! g45n1svt m=1 l=45n w=120n
.ENDS


* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : mux_x1                                       *
* Netlisted  : Tue Nov 25 18:50:48 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764107443711                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764107443711 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764107443711

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764107443712                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764107443712 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764107443712

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_764107443714                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_764107443714 1 2
** N=2 EP=2 FDC=0
.ends M1_NWELL_CDNS_764107443714

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764107443716                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764107443716 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764107443716

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764107443710                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764107443710 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.46017 scb=0.000436376 scc=1.63659e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764107443710

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764107443711                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764107443711 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_764107443711

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv_x1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv_x1 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X0 2 M2_M1_CDNS_764107443716 $T=980 1840 0 0 $X=900 $Y=1710
X1 4 2 1 nmos1v_CDNS_764107443710 $T=640 820 0 0 $X=220 $Y=620
X2 3 2 1 4 pmos1v_CDNS_764107443711 $T=640 2850 0 0 $X=220 $Y=2650
.ends inv_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764107443712                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764107443712 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 3 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.32e-14 AS=2.32e-14 PD=6.1e-07 PS=6.1e-07 fw=1.45e-07 sa=5.5e-07 sb=3.45e-07 sca=23.8155 scb=0.0247027 scc=0.0021592 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764107443712

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764107443714                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764107443714 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=5.55e-07 sb=1.4e-07 sca=4.46017 scb=0.000436376 scc=1.63659e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764107443714

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764107443715                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764107443715 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.92e-14 PD=3.6e-07 PS=5.6e-07 fw=1.2e-07 sa=4.5e-07 sb=2.45e-07 sca=4.46017 scb=0.000436376 scc=1.63659e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764107443715

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764107443716                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764107443716 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.32e-14 PD=5.7e-07 PS=6.1e-07 fw=1.45e-07 sa=7.55e-07 sb=1.4e-07 sca=23.8155 scb=0.0247027 scc=0.0021592 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764107443716

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764107443717                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764107443717 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 3 2 1 5 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.32e-14 AS=2.03e-14 PD=6.1e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=7.55e-07 sca=23.8541 scb=0.0247101 scc=0.0021592 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764107443717

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764107443718                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764107443718 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 3 1 2 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.32e-14 AS=2.32e-14 PD=6.1e-07 PS=6.1e-07 fw=1.45e-07 sa=3.45e-07 sb=5.5e-07 sca=23.8155 scb=0.0247027 scc=0.0021592 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764107443718

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mux_x1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mux_x1 10 1 7 5 4 3
** N=11 EP=6 FDC=12
X0 1 M1_PO_CDNS_764107443711 $T=1310 1360 0 0 $X=1210 $Y=1240
X1 2 M1_PO_CDNS_764107443711 $T=2470 1950 0 90 $X=2350 $Y=1850
X2 2 M2_M1_CDNS_764107443712 $T=1120 1840 0 0 $X=900 $Y=1710
X3 1 M2_M1_CDNS_764107443712 $T=3500 1800 0 180 $X=3280 $Y=1670
X4 3 4 M1_NWELL_CDNS_764107443714 $T=2620 3690 0 90 $X=1900 $Y=3390
X5 5 M2_M1_CDNS_764107443716 $T=400 1860 0 0 $X=320 $Y=1730
X6 1 M2_M1_CDNS_764107443716 $T=1310 1360 0 0 $X=1230 $Y=1230
X7 5 2 3 4 inv_x1 $T=0 0 0 0 $X=0 $Y=0
X8 6 7 3 4 inv_x1 $T=4020 0 0 0 $X=4020 $Y=0
X9 8 2 3 4 pmos1v_CDNS_764107443712 $T=2590 2850 1 180 $X=2140 $Y=2650
X10 6 1 9 4 nmos1v_CDNS_764107443714 $T=1970 820 1 180 $X=1460 $Y=620
X11 6 10 11 4 nmos1v_CDNS_764107443714 $T=2710 820 0 0 $X=2510 $Y=620
X12 4 5 9 nmos1v_CDNS_764107443715 $T=2180 820 1 180 $X=1890 $Y=620
X13 6 5 8 4 3 pmos1v_CDNS_764107443716 $T=2180 2850 1 180 $X=1670 $Y=2650
X14 6 1 8 4 3 pmos1v_CDNS_764107443717 $T=3410 2850 1 180 $X=3080 $Y=2650
X15 8 3 10 4 pmos1v_CDNS_764107443718 $T=3000 2850 1 180 $X=2550 $Y=2650
M0 11 2 4 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.92e-14 PD=3.6e-07 PS=5.6e-07 fw=1.2e-07 sa=4.5e-07 sb=2.45e-07 sca=4.46017 scb=0.000436376 scc=1.63659e-07 $X=2500 $Y=820 $dt=0
M1 2 5 3 3 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=31.4202 scb=0.0358526 scc=0.00253079 $X=640 $Y=2850 $dt=1
M2 7 6 3 3 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=31.9453 scb=0.0366664 scc=0.00259967 $X=4660 $Y=2850 $dt=1
.ends mux_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : buffer_x1                                    *
* Netlisted  : Mon Sep  8 17:57:38 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_757365051520                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_757365051520 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.46017 scb=0.000436376 scc=1.63659e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_757365051520

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv_x1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv_x1 Vin Vout vdd! gnd!
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X0 gnd! Vout Vin nmos1v_CDNS_757365051520 $T=640 820 0 0 $X=220 $Y=620
.ends inv_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: buffer_x1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt buffer_x1 gnd! in out vdd!
** N=5 EP=4 FDC=4
X0 in 2 vdd! gnd! inv_x1 $T=0 0 0 0 $X=0 $Y=0
X1 2 out vdd! gnd! inv_x1 $T=1350 0 0 0 $X=1350 $Y=0
M0 2 in vdd! vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=32.74 scb=0.0369217 scc=0.00282966 $X=640 $Y=2850 $dt=1
M1 out 2 vdd! vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=33.2459 scb=0.0377318 scc=0.00289854 $X=1990 $Y=2850 $dt=1
.ends buffer_x1

************************************************************************
* auCdl Netlist:
* 
* Library Name:  watto
* Top Cell Name: latchsr_x1
* View Name:     schematic
* Netlisted on:  Nov 25 20:33:16 2025
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL vdd!
+        gnd!

*.PIN vdd!
*+    gnd!

************************************************************************
* Library Name: watto
* Cell Name:    latchsr_x1
* View Name:    schematic
************************************************************************

.SUBCKT latchsr_x1 Q Qbar Reset Set
*.PININFO Reset:I Set:I Q:O Qbar:O
MPM3 Q Qbar net12 vdd! g45p1svt m=1 l=45n w=145n
MPM2 net12 Reset vdd! vdd! g45p1svt m=1 l=45n w=145n
MPM1 Qbar Q net4 vdd! g45p1svt m=1 l=45n w=145n
MPM0 net4 Set vdd! vdd! g45p1svt m=1 l=45n w=145n
MNM3 Q Reset gnd! gnd! g45n1svt m=1 l=45n w=120n
MNM2 Q Qbar gnd! gnd! g45n1svt m=1 l=45n w=120n
MNM1 Qbar Q gnd! gnd! g45n1svt m=1 l=45n w=120n
MNM0 Qbar Set gnd! gnd! g45n1svt m=1 l=45n w=120n
.ENDS


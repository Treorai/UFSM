* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : nand_x1                                      *
* Netlisted  : Wed Nov 26 18:03:27 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764191003190                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764191003190 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764191003190

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764191003191                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764191003191 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764191003191

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_764191003192                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_764191003192 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_764191003192

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_764191003193                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_764191003193 1 2
** N=2 EP=2 FDC=0
.ends M1_NWELL_CDNS_764191003193

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764191003190                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764191003190 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 3 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.74923 scb=0.000663449 scc=4.92991e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764191003190

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764191003191                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764191003191 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 2 3 1 5 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=33.2274 scb=0.0325337 scc=0.00341592 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764191003191

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nand_x1                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nand_x1 2 1 3 4 5
** N=6 EP=5 FDC=4
X0 1 M1_PO_CDNS_764191003190 $T=510 1570 0 90 $X=390 $Y=1470
X1 2 M1_PO_CDNS_764191003190 $T=510 2050 0 90 $X=390 $Y=1950
X2 1 M1_PO_CDNS_764191003190 $T=1570 1590 0 90 $X=1450 $Y=1490
X3 1 M1_PO_CDNS_764191003190 $T=1570 2240 0 90 $X=1450 $Y=2140
X4 1 M2_M1_CDNS_764191003191 $T=520 1570 0 90 $X=390 $Y=1490
X5 2 M2_M1_CDNS_764191003191 $T=520 2050 0 90 $X=390 $Y=1970
X6 3 M2_M1_CDNS_764191003191 $T=2820 1930 0 0 $X=2740 $Y=1800
X7 4 M1_PSUB_CDNS_764191003192 $T=1480 330 0 90 $X=620 $Y=190
X8 5 4 M1_NWELL_CDNS_764191003193 $T=1600 3690 0 90 $X=880 $Y=3390
X9 4 6 1 4 nmos1v_CDNS_764191003190 $T=860 940 0 0 $X=440 $Y=740
X10 6 3 2 4 nmos1v_CDNS_764191003190 $T=2260 940 0 0 $X=1840 $Y=740
X11 5 3 2 4 5 pmos1v_CDNS_764191003191 $T=860 2790 0 0 $X=440 $Y=2590
X12 3 5 1 4 5 pmos1v_CDNS_764191003191 $T=2260 2790 0 0 $X=1840 $Y=2590
.ends nand_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : nor_x1                                       *
* Netlisted  : Wed Nov 26 23:24:36 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764210272201                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764210272201 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=4.5148 scb=0.000474692 scc=2.05736e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764210272201

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764210272202                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764210272202 1 2 3
** N=3 EP=3 FDC=1
M0 1 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=4.5148 scb=0.000474692 scc=2.05736e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764210272202

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nor_x1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nor_x1 A B S gnd! vdd!
** N=6 EP=5 FDC=4
X2 gnd! B S nmos1v_CDNS_764210272201 $T=1400 845 1 180 $X=1070 $Y=645
X3 S gnd! A nmos1v_CDNS_764210272202 $T=900 845 0 0 $X=480 $Y=645
M0 3 A S vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=8.7e-15 AS=2.03e-14 PD=4.1e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=2.45e-07 sca=28.9241 scb=0.030769 scc=0.0019811 $X=900 $Y=2865 $dt=1
M1 vdd! B 3 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=8.7e-15 PD=5.7e-07 PS=4.1e-07 fw=1.45e-07 sa=2.45e-07 sb=1.4e-07 sca=29.3918 scb=0.0317277 scc=0.00202057 $X=1110 $Y=2865 $dt=1
.ends nor_x1

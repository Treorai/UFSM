* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : latchsr_x1                                   *
* Netlisted  : Tue Nov 25 20:33:20 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764113596371                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764113596371 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764113596371

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_764113596373                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_764113596373 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_764113596373

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_764113596374                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_764113596374 1 2
** N=2 EP=2 FDC=0
.ends M1_NWELL_CDNS_764113596374

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764113596370                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764113596370 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=4.62022 scb=0.00055476 scc=3.11054e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764113596370

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764113596371                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764113596371 1 2 3
** N=3 EP=3 FDC=1
M0 1 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.62022 scb=0.00055476 scc=3.11054e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764113596371

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764113596372                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764113596372 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_764113596372

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764113596373                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764113596373 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_764113596373

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764113596374                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764113596374 1 2 3
** N=3 EP=3 FDC=1
M0 1 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=4.62022 scb=0.00055476 scc=3.11054e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764113596374

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: latchsr_x1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt latchsr_x1 2 1 6 5 3 4
** N=8 EP=6 FDC=8
X0 1 M1_PO_CDNS_764113596371 $T=1520 2290 0 0 $X=1300 $Y=2170
X1 2 M1_PO_CDNS_764113596371 $T=1850 1540 0 0 $X=1630 $Y=1420
X2 3 M1_PSUB_CDNS_764113596373 $T=2280 300 0 0 $X=1420 $Y=160
X3 4 3 M1_NWELL_CDNS_764113596374 $T=2280 3700 0 0 $X=1380 $Y=3400
X4 3 5 1 nmos1v_CDNS_764113596370 $T=620 890 0 0 $X=200 $Y=690
X5 2 3 1 nmos1v_CDNS_764113596371 $T=2620 890 1 180 $X=2110 $Y=690
X6 2 3 6 nmos1v_CDNS_764113596371 $T=3980 890 0 0 $X=3560 $Y=690
X7 1 2 7 3 4 pmos1v_CDNS_764113596372 $T=1030 2850 0 0 $X=830 $Y=2650
X8 2 1 8 3 4 pmos1v_CDNS_764113596372 $T=2620 2850 1 180 $X=2110 $Y=2650
X9 4 5 7 3 pmos1v_CDNS_764113596373 $T=820 2850 0 0 $X=400 $Y=2650
X10 4 6 8 3 pmos1v_CDNS_764113596373 $T=2830 2850 1 180 $X=2540 $Y=2650
X11 1 3 2 nmos1v_CDNS_764113596374 $T=1120 890 1 180 $X=670 $Y=690
M0 7 5 4 4 g45p1svt L=4.5e-08 W=1.45e-07 AD=8.7e-15 AS=2.03e-14 PD=4.1e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=2.45e-07 sca=28.2191 scb=0.0304148 scc=0.00223692 $X=820 $Y=2850 $dt=1
M1 1 2 7 4 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=8.7e-15 PD=5.7e-07 PS=4.1e-07 fw=1.45e-07 sa=2.45e-07 sb=1.4e-07 sca=26.326 scb=0.0271677 scc=0.00217105 $X=1030 $Y=2850 $dt=1
M2 8 1 2 4 g45p1svt L=4.5e-08 W=1.45e-07 AD=8.7e-15 AS=2.03e-14 PD=4.1e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=2.45e-07 sca=23.8155 scb=0.0247027 scc=0.0021592 $X=2530 $Y=2850 $dt=1
M3 4 6 8 4 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=8.7e-15 PD=5.7e-07 PS=4.1e-07 fw=1.45e-07 sa=2.45e-07 sb=1.4e-07 sca=23.9386 scb=0.0247294 scc=0.0021592 $X=2740 $Y=2850 $dt=1
.ends latchsr_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : xnor_x1                                      *
* Netlisted  : Tue Nov 25 17:06:38 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764101194240                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764101194240 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764101194240

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764101194241                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764101194241 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764101194241

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_764101194242                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_764101194242 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_764101194242

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764101194240                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764101194240 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.46017 scb=0.000436376 scc=1.63659e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764101194240

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764101194241                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764101194241 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_764101194241

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv_x1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv_x1 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X0 1 M2_M1_CDNS_764101194241 $T=980 1840 0 0 $X=900 $Y=1710
X1 4 2 1 4 nmos1v_CDNS_764101194240 $T=640 820 0 0 $X=220 $Y=620
X2 3 1 2 4 3 pmos1v_CDNS_764101194241 $T=640 2850 0 0 $X=220 $Y=2650
.ends inv_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xnor_x1                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xnor_x1 2 3 6 7 9
** N=11 EP=5 FDC=12
X0 1 M1_PO_CDNS_764101194240 $T=2380 1860 0 90 $X=2260 $Y=1760
X1 2 M1_PO_CDNS_764101194240 $T=2640 2320 0 90 $X=2520 $Y=2220
X2 1 M1_PO_CDNS_764101194240 $T=3140 1910 0 90 $X=3020 $Y=1810
X3 2 M1_PO_CDNS_764101194240 $T=4110 1960 0 0 $X=4010 $Y=1840
X4 3 M1_PO_CDNS_764101194240 $T=4390 1420 0 90 $X=4270 $Y=1320
X5 2 M1_PO_CDNS_764101194240 $T=4900 1960 0 0 $X=4800 $Y=1840
X6 1 M1_PO_CDNS_764101194240 $T=4950 2320 0 90 $X=4830 $Y=2220
X7 4 M1_PO_CDNS_764101194240 $T=5730 1430 0 90 $X=5610 $Y=1330
X8 4 M1_PO_CDNS_764101194240 $T=7010 2360 0 90 $X=6890 $Y=2260
X9 2 M2_M1_CDNS_764101194241 $T=2650 2320 0 90 $X=2520 $Y=2240
X10 5 M2_M1_CDNS_764101194241 $T=3630 1930 0 90 $X=3500 $Y=1850
X11 3 M2_M1_CDNS_764101194241 $T=4380 1420 0 90 $X=4250 $Y=1340
X12 4 M2_M1_CDNS_764101194241 $T=5730 1430 0 90 $X=5600 $Y=1350
X13 4 M2_M1_CDNS_764101194241 $T=7010 2360 0 90 $X=6880 $Y=2280
X14 6 M2_M1_CDNS_764101194241 $T=7690 2090 0 90 $X=7560 $Y=2010
X15 5 M2_M1_CDNS_764101194241 $T=7700 1720 0 90 $X=7570 $Y=1640
X16 4 M3_M2_CDNS_764101194242 $T=1180 1830 0 0 $X=1100 $Y=1700
X17 5 M3_M2_CDNS_764101194242 $T=3630 1930 0 90 $X=3500 $Y=1850
X18 4 M3_M2_CDNS_764101194242 $T=5270 1430 0 90 $X=5140 $Y=1350
X19 5 M3_M2_CDNS_764101194242 $T=7700 1720 0 90 $X=7570 $Y=1640
X20 7 1 5 7 nmos1v_CDNS_764101194240 $T=3170 820 0 0 $X=2750 $Y=620
X21 7 3 8 7 nmos1v_CDNS_764101194240 $T=4420 820 0 0 $X=4000 $Y=620
X22 8 4 6 7 nmos1v_CDNS_764101194240 $T=5690 1060 1 0 $X=5270 $Y=620
X23 5 2 6 7 nmos1v_CDNS_764101194240 $T=7050 1060 0 180 $X=6540 $Y=620
X24 9 10 2 7 9 pmos1v_CDNS_764101194241 $T=3240 2850 0 0 $X=2820 $Y=2650
X25 10 6 3 7 9 pmos1v_CDNS_764101194241 $T=4420 2850 0 0 $X=4000 $Y=2650
X26 11 6 1 7 9 pmos1v_CDNS_764101194241 $T=5750 3140 0 180 $X=5240 $Y=2650
X27 11 9 4 7 9 pmos1v_CDNS_764101194241 $T=6960 2850 0 0 $X=6540 $Y=2650
X28 4 2 9 7 inv_x1 $T=0 0 0 0 $X=0 $Y=0
X29 1 3 9 7 inv_x1 $T=1350 0 0 0 $X=1350 $Y=0
M0 4 2 9 9 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=31.4202 scb=0.0358526 scc=0.00253079 $X=640 $Y=2850 $dt=1
M1 1 3 9 9 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=23.8249 scb=0.0247044 scc=0.0021592 $X=1990 $Y=2850 $dt=1
M2 10 2 9 9 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=23.8155 scb=0.0247027 scc=0.0021592 $X=3240 $Y=2850 $dt=1
M3 6 3 10 9 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=23.8155 scb=0.0247027 scc=0.0021592 $X=4420 $Y=2850 $dt=1
M4 11 1 6 9 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=23.8155 scb=0.0247027 scc=0.0021592 $X=5660 $Y=2850 $dt=1
M5 9 4 11 9 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.9072 scb=0.0281197 scc=0.00218359 $X=6960 $Y=2850 $dt=1
.ends xnor_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : tristatebuffer_x1                            *
* Netlisted  : Tue Nov 25 20:16:17 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764112572791                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764112572791 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764112572791

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_764112572795                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_764112572795 1
** N=1 EP=1 FDC=0
.ends M1_NWELL_CDNS_764112572795

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_764112572796                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_764112572796 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_764112572796

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764112572790                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764112572790 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.46017 scb=0.000436376 scc=1.63659e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764112572790

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764112572791                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764112572791 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_764112572791

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv_x1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv_x1 1 2 3 4
** N=4 EP=4 FDC=2
X0 3 M1_NWELL_CDNS_764112572795 $T=670 3700 0 0 $X=130 $Y=3400
X1 4 M1_PSUB_CDNS_764112572796 $T=680 300 0 0 $X=180 $Y=160
X2 4 2 1 nmos1v_CDNS_764112572790 $T=640 820 0 0 $X=220 $Y=620
X3 3 2 1 4 pmos1v_CDNS_764112572791 $T=640 2850 0 0 $X=220 $Y=2650
M0 2 1 3 3 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=31.4202 scb=0.0358526 scc=0.00253079 $X=640 $Y=2850 $dt=1
.ends inv_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764112572792                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764112572792 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 1 g45p1svt L=4.5e-08 W=1.45e-07 AD=8.7e-15 AS=2.03e-14 PD=4.1e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=2.45e-07 sca=26.5414 scb=0.0263556 scc=0.002507 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764112572792

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764112572793                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764112572793 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=8.7e-15 PD=5.7e-07 PS=4.1e-07 fw=1.45e-07 sa=2.45e-07 sb=1.4e-07 sca=27.3953 scb=0.0274124 scc=0.00251189 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764112572793

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764112572794                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764112572794 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=4.46017 scb=0.000436376 scc=1.63659e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764112572794

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764112572795                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764112572795 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=4.46017 scb=0.000436376 scc=1.63659e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764112572795

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: tristatebuffer_x1                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt tristatebuffer_x1 6 5 1 8 4
** N=9 EP=5 FDC=8
X0 1 M1_PO_CDNS_764112572791 $T=1860 2300 0 0 $X=1520 $Y=2180
X1 2 M1_PO_CDNS_764112572791 $T=2810 1420 0 0 $X=2470 $Y=1300
X2 3 M1_PO_CDNS_764112572791 $T=3260 1880 0 0 $X=2920 $Y=1760
X3 4 M1_NWELL_CDNS_764112572795 $T=2980 3700 0 0 $X=2440 $Y=3400
X4 5 M1_PSUB_CDNS_764112572796 $T=3020 300 0 0 $X=2520 $Y=160
X5 5 2 1 nmos1v_CDNS_764112572790 $T=2200 820 0 0 $X=1780 $Y=620
X6 4 2 1 5 pmos1v_CDNS_764112572791 $T=2200 2840 0 0 $X=1780 $Y=2640
X7 6 3 4 5 inv_x1 $T=0 0 0 0 $X=0 $Y=0
X8 4 2 7 5 pmos1v_CDNS_764112572792 $T=3390 2830 0 0 $X=2970 $Y=2630
X9 8 3 7 5 4 pmos1v_CDNS_764112572793 $T=3600 2830 0 0 $X=3400 $Y=2630
X10 8 6 9 5 nmos1v_CDNS_764112572794 $T=3600 820 0 0 $X=3400 $Y=620
X11 5 2 9 nmos1v_CDNS_764112572795 $T=3390 820 0 0 $X=2970 $Y=620
M0 2 1 4 4 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=24.5515 scb=0.0251693 scc=0.00232652 $X=2200 $Y=2840 $dt=1
.ends tristatebuffer_x1

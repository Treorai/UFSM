* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : 4_bit_full_adder_x1                          *
* Netlisted  : Mon Dec  1 23:41:38 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764643294310                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764643294310 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 3 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.74923 scb=0.000663449 scc=4.92991e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764643294310

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nand_x1                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nand_x1 B A gnd! vdd! S
*.DEVICECLIMB
** N=6 EP=5 FDC=2
X9 gnd! 6 B gnd! nmos1v_CDNS_764643294310 $T=860 940 0 0 $X=440 $Y=740
X10 6 S A gnd! nmos1v_CDNS_764643294310 $T=2260 940 0 0 $X=1840 $Y=740
.ends nand_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 1_bit_full_adder_x1                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 1_bit_full_adder_x1 A B gnd! vdd! CarryIn CarryOut S
** N=23 EP=7 FDC=36
X17 B A gnd! vdd! 8 nand_x1 $T=0 0 0 0 $X=0 $Y=0
X18 B 8 gnd! vdd! 12 nand_x1 $T=3210 0 0 0 $X=3210 $Y=0
X19 12 9 gnd! vdd! 10 nand_x1 $T=6420 0 0 0 $X=6420 $Y=0
X20 8 A gnd! vdd! 9 nand_x1 $T=9630 0 0 0 $X=9630 $Y=0
X21 CarryIn 10 gnd! vdd! 13 nand_x1 $T=12840 0 0 0 $X=12840 $Y=0
X22 CarryIn 13 gnd! vdd! 11 nand_x1 $T=16050 0 0 0 $X=16050 $Y=0
X23 8 13 gnd! vdd! CarryOut nand_x1 $T=19260 0 0 0 $X=19260 $Y=0
X24 13 10 gnd! vdd! 14 nand_x1 $T=22470 0 0 0 $X=22470 $Y=0
X25 11 14 gnd! vdd! S nand_x1 $T=25680 0 0 0 $X=25680 $Y=0
M0 8 A vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=30.5075 scb=0.0298234 scc=0.00339941 $X=860 $Y=2790 $dt=1
M1 vdd! B 8 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=2260 $Y=2790 $dt=1
M2 12 8 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=4070 $Y=2790 $dt=1
M3 vdd! B 12 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=5470 $Y=2790 $dt=1
M4 10 9 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=7280 $Y=2790 $dt=1
M5 vdd! 12 10 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=8680 $Y=2790 $dt=1
M6 9 A vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=10490 $Y=2790 $dt=1
M7 vdd! 8 9 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=11890 $Y=2790 $dt=1
M8 13 10 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=13700 $Y=2790 $dt=1
M9 vdd! CarryIn 13 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=15100 $Y=2790 $dt=1
M10 11 13 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=16910 $Y=2790 $dt=1
M11 vdd! CarryIn 11 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=18310 $Y=2790 $dt=1
M12 CarryOut 13 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=20120 $Y=2790 $dt=1
M13 vdd! 8 CarryOut vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=21520 $Y=2790 $dt=1
M14 14 10 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=23330 $Y=2790 $dt=1
M15 vdd! 13 14 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=24730 $Y=2790 $dt=1
M16 S 14 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.5685 scb=0.0249349 scc=0.00334489 $X=26540 $Y=2790 $dt=1
M17 vdd! 11 S vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=30.5075 scb=0.0298234 scc=0.00339941 $X=27940 $Y=2790 $dt=1
.ends 1_bit_full_adder_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 4_bit_full_adder_x1                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 4_bit_full_adder_x1 A0 A1 A2 A3 B0 B1 B2 B3 CarryIn CarryOut
+ S0 S1 S2 S3 gnd! vdd!
** N=83 EP=16 FDC=144
X14 A0 B0 gnd! vdd! CarryIn 6 S0 1_bit_full_adder_x1 $T=0 0 0 0 $X=0 $Y=0
X15 A1 B1 gnd! vdd! 6 10 S1 1_bit_full_adder_x1 $T=0 8000 1 0 $X=0 $Y=4000
X16 A2 B2 gnd! vdd! 10 14 S2 1_bit_full_adder_x1 $T=0 8000 0 0 $X=0 $Y=8000
X17 A3 B3 gnd! vdd! 14 CarryOut S3 1_bit_full_adder_x1 $T=0 16000 1 0 $X=0 $Y=12000
.ends 4_bit_full_adder_x1

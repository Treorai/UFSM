* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : nand_x1                                      *
* Netlisted  : Wed Nov 26 18:03:27 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764191003190                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764191003190 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 3 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.74923 scb=0.000663449 scc=4.92991e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764191003190

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764191003191                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764191003191 1 2 3 5
** N=5 EP=4 FDC=1
M0 2 3 1 5 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=33.2274 scb=0.0325337 scc=0.00341592 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764191003191

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nand_x1                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nand_x1 A B S gnd! vdd!
** N=6 EP=5 FDC=4
X9 gnd! 6 B gnd! nmos1v_CDNS_764191003190 $T=860 940 0 0 $X=440 $Y=740
X10 6 S A gnd! nmos1v_CDNS_764191003190 $T=2260 940 0 0 $X=1840 $Y=740
X11 vdd! S A vdd! pmos1v_CDNS_764191003191 $T=860 2790 0 0 $X=440 $Y=2590
X12 S vdd! B vdd! pmos1v_CDNS_764191003191 $T=2260 2790 0 0 $X=1840 $Y=2590
.ends nand_x1

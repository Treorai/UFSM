library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mod is
end mod;

architecture Behavioral of mod is

begin


end Behavioral;


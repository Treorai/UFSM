* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : switch_x1                                    *
* Netlisted  : Tue Nov 25 17:40:56 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764103252230                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764103252230 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764103252230

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764103252231                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764103252231 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764103252231

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764103252230                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764103252230 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_764103252230

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764103252231                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764103252231 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 3 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.46017 scb=0.000436376 scc=1.63659e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764103252231

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv_x1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv_x1 1 2 3 4
** N=4 EP=4 FDC=2
X0 2 M2_M1_CDNS_764103252231 $T=980 1840 0 0 $X=900 $Y=1710
X1 4 2 1 3 4 pmos1v_CDNS_764103252230 $T=640 2850 0 0 $X=220 $Y=2650
X2 3 2 1 3 nmos1v_CDNS_764103252231 $T=640 820 0 0 $X=220 $Y=620
M0 2 1 4 4 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=31.4202 scb=0.0358526 scc=0.00253079 $X=640 $Y=2850 $dt=1
.ends inv_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: switch_x1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt switch_x1 2 3 4 5 6
** N=6 EP=5 FDC=4
X0 1 M1_PO_CDNS_764103252230 $T=1020 1860 0 90 $X=900 $Y=1760
X1 2 M1_PO_CDNS_764103252230 $T=1320 1420 0 90 $X=1200 $Y=1320
X2 2 M2_M1_CDNS_764103252231 $T=1330 1420 0 90 $X=1200 $Y=1340
X3 3 M2_M1_CDNS_764103252231 $T=1820 2290 0 0 $X=1740 $Y=2160
X4 4 M2_M1_CDNS_764103252231 $T=1840 950 0 0 $X=1760 $Y=820
X5 4 M2_M1_CDNS_764103252231 $T=2510 2240 0 0 $X=2430 $Y=2110
X6 3 4 1 5 6 pmos1v_CDNS_764103252230 $T=2000 2850 0 0 $X=1580 $Y=2650
X7 4 3 2 5 nmos1v_CDNS_764103252231 $T=2000 820 0 0 $X=1580 $Y=620
X8 2 1 5 6 inv_x1 $T=0 0 0 0 $X=0 $Y=0
M0 4 1 3 6 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=29.9008 scb=0.0333585 scc=0.00236277 $X=2000 $Y=2850 $dt=1
.ends switch_x1

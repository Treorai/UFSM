* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : flipflopD_barless_x1                         *
* Netlisted  : Sat Nov 29 19:17:02 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764454616470                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764454616470 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.92313 scb=0.000827672 scc=8.57018e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764454616470

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764454616472                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764454616472 1 2 3
** N=4 EP=3 FDC=1
M0 1 2 3 3 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.32e-14 PD=5.7e-07 PS=6.1e-07 fw=1.45e-07 sa=3.45e-07 sb=1.4e-07 sca=22.508 scb=0.0238066 scc=0.00185903 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764454616472

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764454616473                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764454616473 1 2 3
** N=4 EP=3 FDC=1
M0 2 3 1 1 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.32e-14 AS=2.03e-14 PD=6.1e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=3.45e-07 sca=22.508 scb=0.0238066 scc=0.00185903 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764454616473

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764454616474                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764454616474 1 2 3 5
** N=5 EP=4 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.32e-14 PD=5.7e-07 PS=6.1e-07 fw=1.45e-07 sa=3.45e-07 sb=1.4e-07 sca=22.508 scb=0.0238066 scc=0.00185903 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764454616474

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764454616475                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764454616475 1 2 3
** N=4 EP=3 FDC=1
M0 2 3 1 1 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.32e-14 PD=5.7e-07 PS=6.1e-07 fw=1.45e-07 sa=3.45e-07 sb=1.4e-07 sca=22.508 scb=0.0238066 scc=0.00185903 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764454616475

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764454616476                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764454616476 1 2 3
** N=3 EP=3 FDC=1
M0 1 2 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=4.92313 scb=0.000827672 scc=8.57018e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764454616476

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764454616477                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764454616477 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=4.92313 scb=0.000827672 scc=8.57018e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764454616477

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: flipflopD_barless_x1                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt flipflopD_barless_x1 D Q clk gnd! vdd!
** N=10 EP=5 FDC=12
X18 gnd! 5 3 gnd! nmos1v_CDNS_764454616470 $T=720 1000 0 0 $X=300 $Y=800
X19 gnd! 3 7 gnd! nmos1v_CDNS_764454616470 $T=2500 1000 0 0 $X=2080 $Y=800
X20 5 clk D gnd! nmos1v_CDNS_764454616470 $T=4380 1000 0 0 $X=3960 $Y=800
X21 Q clk 6 gnd! nmos1v_CDNS_764454616470 $T=7790 1000 0 0 $X=7370 $Y=800
X24 Q 10 vdd! pmos1v_CDNS_764454616472 $T=6390 2870 0 0 $X=6150 $Y=2670
X25 vdd! 7 3 pmos1v_CDNS_764454616473 $T=2500 2870 0 0 $X=2080 $Y=2670
X26 6 clk 7 vdd! pmos1v_CDNS_764454616474 $T=2910 2870 0 0 $X=2670 $Y=2670
X27 vdd! 10 6 pmos1v_CDNS_764454616475 $T=6070 2870 1 180 $X=5560 $Y=2670
X28 Q 10 gnd! nmos1v_CDNS_764454616476 $T=6390 1000 0 0 $X=6150 $Y=800
X29 gnd! 10 6 nmos1v_CDNS_764454616477 $T=6070 1000 1 180 $X=5560 $Y=800
M0 3 5 vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=28.4097 scb=0.0321484 scc=0.00204568 $X=720 $Y=2870 $dt=1
M1 7 clk 5 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=22.508 scb=0.0238066 scc=0.00185903 $X=4380 $Y=2870 $dt=1
.ends flipflopD_barless_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : xnor_x1                                      *
* Netlisted  : Tue Nov 25 17:06:38 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764101194240                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764101194240 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.46017 scb=0.000436376 scc=1.63659e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764101194240

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv_x1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv_x1 Vout Vin vdd! gnd!
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X1 gnd! Vin Vout gnd! nmos1v_CDNS_764101194240 $T=640 820 0 0 $X=220 $Y=620
.ends inv_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: xnor_x1                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt xnor_x1 A B S gnd! vdd!
** N=11 EP=5 FDC=12
X20 gnd! 1 5 gnd! nmos1v_CDNS_764101194240 $T=3170 820 0 0 $X=2750 $Y=620
X21 gnd! B 8 gnd! nmos1v_CDNS_764101194240 $T=4420 820 0 0 $X=4000 $Y=620
X22 8 4 S gnd! nmos1v_CDNS_764101194240 $T=5690 1060 1 0 $X=5270 $Y=620
X23 5 A S gnd! nmos1v_CDNS_764101194240 $T=7050 1060 0 180 $X=6540 $Y=620
X28 4 A vdd! gnd! inv_x1 $T=0 0 0 0 $X=0 $Y=0
X29 1 B vdd! gnd! inv_x1 $T=1350 0 0 0 $X=1350 $Y=0
M0 4 A vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=31.4202 scb=0.0358526 scc=0.00253079 $X=640 $Y=2850 $dt=1
M1 1 B vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=23.8249 scb=0.0247044 scc=0.0021592 $X=1990 $Y=2850 $dt=1
M2 10 A vdd! vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=23.8155 scb=0.0247027 scc=0.0021592 $X=3240 $Y=2850 $dt=1
M3 S B 10 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=23.8155 scb=0.0247027 scc=0.0021592 $X=4420 $Y=2850 $dt=1
M4 11 1 S vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=23.8155 scb=0.0247027 scc=0.0021592 $X=5660 $Y=2850 $dt=1
M5 vdd! 4 11 vdd! g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=26.9072 scb=0.0281197 scc=0.00218359 $X=6960 $Y=2850 $dt=1
.ends xnor_x1

************************************************************************
* auCdl Netlist:
* 
* Library Name:  watto
* Top Cell Name: buffer_x2
* View Name:     schematic
* Netlisted on:  Nov 25 18:37:23 2025
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL vdd!
+        gnd!

*.PIN vdd!
*+    gnd!

************************************************************************
* Library Name: watto
* Cell Name:    inv_x2
* View Name:    schematic
************************************************************************

.SUBCKT inv_x2 Vin Vout
*.PININFO Vin:I Vout:O
MNM0 Vout Vin gnd! gnd! g45n1svt m=1 l=45n w=240n
MPM0 Vout Vin vdd! vdd! g45p1svt m=1 l=45n w=290n
.ENDS

************************************************************************
* Library Name: watto
* Cell Name:    buffer_x2
* View Name:    schematic
************************************************************************

.SUBCKT buffer_x2 in out
*.PININFO in:I out:O
XI2 in net2 / inv_x2
XI3 net2 out / inv_x2
.ENDS


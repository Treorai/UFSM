* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : tristateinv_x1                               *
* Netlisted  : Tue Nov 25 19:42:28 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764110544150                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764110544150 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=4.3585 scb=0.000370956 scc=1.03875e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764110544150

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764110544151                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764110544151 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.46017 scb=0.000436376 scc=1.63659e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764110544151

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764110544152                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764110544152 1 2 3
** N=4 EP=3 FDC=1
M0 2 3 1 1 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=2.03e-14 PD=5.7e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=1.4e-07 sca=31.4202 scb=0.0358526 scc=0.00253079 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764110544152

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv_x1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv_x1 Vin Vout vdd! gnd!
** N=4 EP=4 FDC=2
X2 gnd! Vout Vin nmos1v_CDNS_764110544151 $T=640 820 0 0 $X=220 $Y=620
X3 vdd! Vout Vin pmos1v_CDNS_764110544152 $T=640 2850 0 0 $X=220 $Y=2650
.ends inv_x1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764110544153                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764110544153 1 2 3 5
** N=5 EP=4 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.45e-07 AD=2.03e-14 AS=8.7e-15 PD=5.7e-07 PS=4.1e-07 fw=1.45e-07 sa=2.45e-07 sb=1.4e-07 sca=28.3455 scb=0.0306395 scc=0.00224409 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764110544153

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764110544154                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764110544154 1 2 3
** N=4 EP=3 FDC=1
M0 3 2 1 1 g45p1svt L=4.5e-08 W=1.45e-07 AD=8.7e-15 AS=2.03e-14 PD=4.1e-07 PS=5.7e-07 fw=1.45e-07 sa=1.4e-07 sb=2.45e-07 sca=26.3915 scb=0.0272714 scc=0.00217217 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764110544154

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764110544155                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764110544155 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=4.3585 scb=0.000370956 scc=1.03875e-07 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764110544155

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: tristateinv_x1                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt tristateinv_x1 Vin Vout en gnd! vdd!
** N=8 EP=5 FDC=6
X2 Vout Vin 5 gnd! nmos1v_CDNS_764110544150 $T=2230 770 0 0 $X=2030 $Y=570
X3 en 7 vdd! gnd! inv_x1 $T=0 0 0 0 $X=0 $Y=0
X4 Vout Vin 8 vdd! pmos1v_CDNS_764110544153 $T=2230 2850 0 0 $X=2030 $Y=2650
X5 vdd! 7 8 pmos1v_CDNS_764110544154 $T=2020 2850 0 0 $X=1600 $Y=2650
X6 gnd! en 5 nmos1v_CDNS_764110544155 $T=2020 770 0 0 $X=1600 $Y=570
.ends tristateinv_x1

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity a3 is
    Port ( a, b, c, d : in  STD_LOGIC;
           s : out  STD_LOGIC);
end a3;

architecture Behavioral of a3 is

begin


end Behavioral;

